
.subckt 000006_output
m0 net1 net2 gnd gnd nmos4
r1 net0 net1 r
.ends
