
.subckt 000146_output
m0 net3 net3 net0 net0 pmos4
m1 net2 net5 net6 net6 nmos4
m2 net10 net12 gnd gnd nmos4
m3 net8 net11 net10 net10 nmos4
m4 net2 net1 net0 net0 pmos4
m5 net6 net9 net10 net10 nmos4
m6 net3 net7 net8 net8 nmos4
r7 net6 net8 r
.ends
