
.subckt 000164_output
m0 net1 net3 gnd gnd nmos4
r1 net0 net1 r
m2 net2 net4 gnd gnd nmos4
r3 net0 net2 r
.ends
