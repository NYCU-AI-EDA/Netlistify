
.subckt 000157_output
m0 net2 net5 net6 net6 nmos4
m1 net3 net4 net6 net6 nmos4
r2 net0 net2 r
r3 net7 net7 r
r4 net1 net3 r
.ends
