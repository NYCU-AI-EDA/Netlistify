
.subckt 000149_output
m0 net9 net10 gnd gnd nmos4
m1 net2 net1 net0 net0 pmos4
m2 net5 net3 net0 net0 pmos4
m3 net3 net8 net9 net9 nmos4
m4 net6 net7 net9 net9 nmos4
r5 net2 net6 r
r6 net5 net3 r
.ends
