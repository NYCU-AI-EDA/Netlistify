
.subckt 000174_output
m0 net2 net1 gnd gnd nmos4
m1 net0 net1 net2 net2 nmos4
.ends
