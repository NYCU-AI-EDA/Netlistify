
.subckt 000010_output
m0 net1 net2 gnd gnd nmos4
r1 net0 net1 r
r2 net1 gnd r
.ends
