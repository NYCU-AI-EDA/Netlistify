
.subckt 000352_output
m0 net0 net2 net4 net4 nmos4
r1 net5 net7 r
q2 net1 net4 net5 npn
r3 net4 net6 r
r4 net0 net1 r
.ends
