
.subckt 000085_output
m0 net2 net1 net0 net0 pmos4
m1 net1 net3 net5 net5 nmos4
r2 net5 net6 r
r3 net2 gnd r
r4 net5 gnd r
r5 net0 net1 r
.ends
