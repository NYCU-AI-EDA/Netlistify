
.subckt 000356_output
m0 net6 net3 net3 net3 pmos4
m1 net3 net2 net0 net0 pmos4
m2 net4 net6 net7 net7 nmos4
m3 net4 net5 net3 net3 pmos4
m4 net6 net6 net7 net7 nmos4
.ends
