
.subckt 000180_output
v0 net3 gnd v
m1 net2 net4 gnd gnd nmos4
m2 net0 net1 net2 net2 nmos4
.ends
