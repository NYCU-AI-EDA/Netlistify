
.subckt 000348_output
m0 net4 net2 net0 net0 pmos4
m1 net4 net4 net5 net5 nmos4
m2 net4 net1 net0 net0 pmos4
.ends
