
.subckt 000396_output
v0 net3 gnd v
v1 gnd net4 v
i2 net8 net10 i
q3 net2 net4 net6 npn
r4 net5 net8 r
r5 net0 net2 r
r6 net6 net8 r
q7 net1 net3 net5 npn
r8 net0 net1 r
.ends
