
.subckt 000139_output
m0 net2 net2 net0 net0 pmos4
m1 net2 net6 net7 net7 nmos4
m2 net3 net5 net8 net8 nmos4
m3 net8 net9 gnd gnd nmos4
m4 net3 net2 net1 net1 pmos4
.ends
