
.subckt 000053_output
m0 net7 net3 net0 net0 pmos4
m1 net2 net1 net0 net0 pmos4
m2 net4 net2 net0 net0 pmos4
m3 net3 net1 net0 net0 pmos4
m4 net7 net9 gnd gnd nmos4
i5 net6 gnd i
m6 net4 net9 gnd gnd nmos4
m7 net3 net5 net6 net6 nmos4
m8 net2 net8 net6 net6 nmos4
.ends
