
.subckt 000110_output
m0 net3 net1 net0 net0 pmos4
m1 net5 net7 gnd gnd nmos4
m2 net3 net4 net5 net5 nmos4
r3 net1 net2 r
r4 net7 net5 r
c5 net1 net5 c
c8 gnd net7 c
.ends
