
.subckt 000280_output
q0 net3 net5 net5 npn
r1 net2 net7 r
r2 net1 net2 r
r3 net0 net3 r
r4 net5 net7 r
r5 net4 net8 r
c7 net3 net4 c
c8 net6 net8 c
c9 net2 net2 c
.ends
