
.subckt 000324_output
r0 net0 net2 r
r1 net0 net1 r
i2 net8 net9 i
q3 net1 net6 net8 npn
q4 net5 net7 net8 npn
.ends
