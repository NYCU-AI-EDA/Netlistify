
.subckt 000121_output
m0 net1 net3 net0 net0 pmos4
m1 net1 net3 gnd gnd nmos4
r2 net2 net3 r
.ends
