
.subckt 000096_output
m0 net2 net1 gnd gnd nmos4
r1 net1 net2 r
r2 net0 net2 r
.ends
