
.subckt 000154_output
m0 net5 net6 gnd gnd nmos4
m1 net1 net3 net4 net4 nmos4
m2 net2 net5 net5 net5 nmos4
r3 net0 net1 r
r4 net0 net2 r
.ends
