
.subckt 000220_output
i0 net0 net1 i
m1 net4 net4 net2 net2 pmos4
i2 net4 gnd i
m3 net1 net8 net7 net7 nmos4
m4 net2 net2 net0 net0 pmos4
m5 net5 net4 net3 net3 pmos4
m6 net3 net2 net0 net0 pmos4
m7 net7 net7 gnd gnd nmos4
m8 net9 net10 gnd gnd nmos4
m9 net5 net8 net9 net9 nmos4
.ends
