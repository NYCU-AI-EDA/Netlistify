
.subckt 000124_output
m0 net2 net3 net5 net5 nmos4
m1 net1 net3 gnd gnd nmos4
r2 net0 net1 r
r3 net0 net2 r
r4 net5 gnd r
.ends
