
.subckt 000388_output
v0 net4 gnd v
m1 net2 net1 net0 net0 pmos4
v2 net6 gnd v
m3 net1 net1 net0 net0 pmos4
m4 net2 net6 net5 net5 nmos4
m5 net1 net4 net5 net5 nmos4
i6 net5 net9 i
.ends
