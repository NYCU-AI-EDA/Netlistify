
.subckt 000092_output
m0 net1 net2 net3 net3 nmos4
r1 net0 net1 r
r2 net3 gnd r
.ends
