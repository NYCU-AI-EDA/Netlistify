
.subckt 000117_output
m0 net1 net6 net6 net6 nmos4
m1 net2 net6 net8 net8 nmos4
r2 net0 net1 r
r3 net0 net2 r
c5 net7 gnd c
r6 net7 gnd r
c8 net3 net3 c
c11 net2 gnd c
.ends
