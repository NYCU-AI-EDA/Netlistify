
.subckt 000359_output
m0 net7 gnd net3 net3 pmos4
m1 net5 gnd net3 net3 pmos4
m2 net7 net7 gnd gnd nmos4
m3 net5 net7 gnd gnd nmos4
m4 net2 net8 gnd gnd nmos4
r5 net0 net3 r
r6 gnd net2 r
.ends
