
.subckt 000128_output
m0 net2 net1 gnd gnd nmos4
m1 net1 net1 gnd gnd nmos4
r2 net0 net1 r
r3 net0 net2 r
.ends
