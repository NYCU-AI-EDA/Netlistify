
.subckt 000183_output
v0 net1 gnd v
m1 net1 net2 gnd gnd nmos4
r2 net0 net1 r
.ends
