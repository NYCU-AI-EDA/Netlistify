
.subckt 000381_output
m0 net3 net1 net0 net0 pmos4
m1 net8 net1 net0 net0 pmos4
m2 net5 net4 net3 net3 pmos4
m3 net6 net7 net3 net3 pmos4
m4 net6 net5 net10 net10 nmos4
m5 net1 net1 net0 net0 pmos4
m6 net11 net6 net10 net10 nmos4
i7 net1 net10 i
m8 net5 net5 net10 net10 nmos4
c10 net6 net8 c
.ends
