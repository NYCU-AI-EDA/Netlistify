
.subckt 000340_output
m0 net2 net1 net0 net0 pmos4
m1 net3 net1 net0 net0 pmos4
m2 net3 net4 net6 net6 nmos4
m3 net2 net5 net6 net6 nmos4
.ends
