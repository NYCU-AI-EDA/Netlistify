
.subckt 000270_output
i0 net0 net1 i
m1 net3 net2 net4 net4 nmos4
m2 net4 net4 gnd gnd nmos4
.ends
