
.subckt 000311_output
i0 gnd net0 i
q1 net1 net1 net1 npn
r2 net1 net1 r
.ends
