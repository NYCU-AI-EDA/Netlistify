
.subckt 000325_output
r0 net0 net1 r
m1 net1 net2 gnd gnd nmos4
.ends
