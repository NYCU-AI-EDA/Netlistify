
.subckt 000076_output
m0 net7 net3 gnd gnd nmos4
r1 net6 gnd r
r2 net0 net3 r
m3 net3 net4 net6 net6 nmos4
r4 net1 net7 r
r5 net6 net7 r
r7 net0 net7 r
.ends
