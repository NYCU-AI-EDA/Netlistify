
.subckt 000101_output
m0 net4 net5 net1 net1 pmos4
m1 net1 net2 gnd gnd nmos4
r2 net0 net1 r
r3 net4 net4 r
.ends
