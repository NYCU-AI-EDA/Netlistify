
.subckt 000039_output
i0 net0 net2 i
i1 net1 gnd i
c2 net2 net2 c
c5 net1 net2 c
.ends
