
.subckt 000189_output
m0 net2 net1 net0 net0 pmos4
m1 net2 net3 gnd gnd nmos4
r2 net0 net2 r
.ends
