
.subckt 000397_output
i0 net3 gnd i
q1 net0 net1 net2 npn
q2 net0 net2 net4 npn
.ends
