
.subckt 000316_output
v0 net4 gnd v
v1 net3 gnd v
i2 net8 net9 i
q3 net2 net4 net6 npn
r4 net0 net2 r
q5 net1 net3 net5 npn
r6 net6 net8 r
r7 net5 net8 r
r8 net1 net1 r
.ends
