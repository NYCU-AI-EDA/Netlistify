
.subckt 000058_output
m0 net1 net1 net0 net0 pmos4
m1 net5 net5 net0 net0 pmos4
m2 net2 net1 net0 net0 pmos4
m3 net5 net5 net0 net0 pmos4
i4 net14 gnd i
m5 net4 net8 net8 net8 nmos4
m6 net5 net12 net9 net9 nmos4
i7 net9 gnd i
m8 net5 net12 net13 net13 nmos4
m9 net2 net8 net9 net9 nmos4
c10 gnd gnd c
c13 net6 gnd c
.ends
