
.subckt 000018_output
i0 net7 gnd i
m1 net4 net2 net0 net0 pmos4
m2 net3 net1 net0 net0 pmos4
v3 net5 net6 v
m4 net3 net6 net7 net7 nmos4
m5 net4 net5 net7 net7 nmos4
.ends
