
.subckt 000248_output
m0 net4 net1 net11 net11 nmos4
m1 net4 net1 net0 net0 pmos4
m2 net9 net10 net11 net11 nmos4
m3 net6 net5 net12 net12 nmos4
m4 net1 net3 net0 net0 pmos4
m5 net5 net8 net9 net9 nmos4
m6 net6 net5 net0 net0 pmos4
m7 net1 net7 net9 net9 nmos4
m8 net5 net3 net0 net0 pmos4
.ends
