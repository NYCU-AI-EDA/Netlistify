
.subckt 000001_output
q0 gnd gnd net9 pnp
q1 gnd gnd net8 pnp
q2 gnd gnd net6 pnp
m3 net3 net3 net0 net0 pmos4
m4 net1 net1 net6 net6 nmos4
m5 net3 net1 net7 net7 nmos4
m6 net5 net4 net0 net0 pmos4
m7 net1 net2 net0 net0 pmos4
r8 net5 net9 r
r9 net7 net8 r
.ends
