
.subckt 000287_output
v0 net2 net4 v
v1 net5 net6 v
v2 net4 net5 v
v3 net6 gnd v
q4 net1 net2 gnd npn
r5 net0 net1 r
c6 net1 gnd c
.ends
