
.subckt 000214_output
v0 net2 gnd v
m1 net0 net1 net2 net2 nmos4
r2 net0 net1 r
r3 net1 net2 r
.ends
