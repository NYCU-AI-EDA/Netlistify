
.subckt 000026_output
m0 net1 net2 net0 net0 pmos4
m1 net4 net3 net0 net0 pmos4
m2 net1 net5 net8 net8 nmos4
m3 net8 net12 gnd gnd nmos4
m4 net4 net7 net8 net8 nmos4
c5 net1 net12 c
c7 net12 net4 c
.ends
