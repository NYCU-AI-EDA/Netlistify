
.subckt 000230_output
m0 net1 net1 net0 net0 pmos4
m1 net2 net3 gnd gnd nmos4
m2 net2 net1 net0 net0 pmos4
r3 net1 gnd r
.ends
