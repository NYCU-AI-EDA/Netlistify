
.subckt 000222_output
i0 net0 net1 i
i1 net0 net2 i
i2 net4 net6 i
m3 net1 net3 net4 net4 nmos4
m4 net2 net5 net4 net4 nmos4
c5 net1 net2 c
.ends
