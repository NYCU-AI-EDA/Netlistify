
.subckt 000198_output
m0 net2 net4 gnd gnd nmos4
m1 net1 net3 net2 net2 nmos4
r2 net0 net1 r
.ends
