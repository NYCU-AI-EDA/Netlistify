
.subckt 000243_output
m0 net3 net3 net0 net0 pmos4
m1 net1 net4 net0 net0 pmos4
m2 net2 net1 net0 net0 pmos4
m3 net4 net3 net0 net0 pmos4
m4 net4 net10 net7 net7 nmos4
m5 net2 net1 net13 net13 nmos4
m6 net5 net2 net0 net0 pmos4
m7 net3 net6 net7 net7 nmos4
m8 net1 net12 net13 net13 nmos4
c9 net5 gnd c
m10 net7 net12 net13 net13 nmos4
m11 net5 net2 net14 net14 nmos4
.ends
