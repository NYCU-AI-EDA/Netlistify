
.subckt 000332_output
q0 net4 net2 net0 pnp
r1 net1 net2 r
r2 net4 gnd r
q3 net2 net4 gnd npn
c6 net3 net4 c
.ends
