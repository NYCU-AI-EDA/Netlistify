
.subckt 000236_output
q0 gnd gnd net2 pnp
r1 net0 net2 r
.ends
