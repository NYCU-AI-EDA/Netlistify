
.subckt 000250_output
i0 net0 net5 i
m1 net2 net2 net0 net0 pmos4
m2 net5 net5 net15 net15 nmos4
m3 net3 net12 net9 net9 nmos4
m4 net4 net1 net0 net0 pmos4
m5 net8 net5 net15 net15 nmos4
m6 net2 net7 net8 net8 nmos4
m7 net3 net2 net0 net0 pmos4
m8 net4 net14 net15 net15 nmos4
m9 net10 net14 net16 net16 nmos4
q10 net0 net6 net10 npn
q11 net0 net4 net6 npn
.ends
