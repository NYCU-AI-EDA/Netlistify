
.subckt 000379_output
m0 net12 net8 net3 net3 pmos4
m1 net3 net4 net0 net0 pmos4
m2 net6 net6 net1 net1 pmos4
m3 net2 net1 net0 net0 pmos4
m4 net1 net1 net0 net0 pmos4
m5 net12 net12 net13 net13 nmos4
m6 net7 net6 net2 net2 pmos4
m7 net11 net10 net13 net13 nmos4
m8 net7 net10 net11 net11 nmos4
i9 net6 net13 i
.ends
