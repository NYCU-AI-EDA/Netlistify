
.subckt 000032_output
m0 net1 net1 net0 net0 pmos4
m1 net4 net1 net0 net0 pmos4
m2 net1 net4 net5 net5 nmos4
m3 net2 net1 net4 net4 nmos4
m4 net4 net4 gnd gnd nmos4
r5 net5 gnd r
.ends
